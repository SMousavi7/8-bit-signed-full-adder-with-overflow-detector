include "fullAdder.v";

module full_Adder_tb();
	reg [7:0]a;
	reg [7:0]b;
	reg Cin;
	wire [7:0]sum;
	wire Cout;

	full_Adder s(sum, Cout, a, b, Cin);
	initial begin
	a = 12;
	b = 17;
	Cin = 0;
	#50;
	a = 16;
	b  = 10;
	Cin = 1;
	#50;
	a = 54;
	b = 21;
	Cin = 0;
	#50;
	a = 127;
	b = 0;
	Cin = 1;
	#50;
	a = 0;
	b = 0; 
	Cin = 1;
	#50;
	a = 127;
	b = -128; 
	Cin = 0;
	#50;
	a = -128;
	b = -128; 
	Cin = 1;
	#50;
	a = 77;
	b = -77; 
	Cin = 1;
	#50;
	a = 45;
	b = 21; 
	Cin = 1;
	#50;
	a = 100;
	b = 97; 
	Cin = 1;
	#50;
	a = -128;
	b = -128; 
	Cin = 0;
	#50;
	a = 100;
	b = -70;
	Cin = 1;
	#50;
	a = -100;
	b = 70;
	Cin = 0;
	#50;
	a = 54;
	b = 91;
	Cin = 1;
	#50;
	a = -54;
	b = -91;
	Cin = 1;
	#50;
	a = -38;	
	b = -107;	
	Cin = 0;
	#50;
	a = 43;
	b = 93;	
	Cin = 1;
	#50;
	end
endmodule
